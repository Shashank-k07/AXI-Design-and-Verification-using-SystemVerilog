`include"axi_tx.sv"
`include"axi_interface.sv"
`include"common.sv"
`include"axi_gen.sv"
`include"axi_bfm.sv"
`include"axi_slave_bfm.sv"
`include"axi_monitor.sv"
`include"axi_scoreboard.sv"
`include"axi_env.sv"
`include"axi_top.sv"
